{"reason": "DDH_ALIVE", "logger_mac": "", "logger_sn": "", "project": "kaz", "vessel": "joaquim", "ddh_commit": "43830", "utc_time": 1683509450, "local_time": 1683495050, "box_sn": "9999999", "hw_uptime": " 21:30:50 up 2 days,  1:52,  1 user,  load average: 0.22, 0.35, 0.55\n", "gps_position": "+38.000000,-83.000000", "platform": "dev", "msg_ver": 1, "data": ""}